entity cla4b is
port();
end cla4b;

architecture cla of cla4b is
begin

end cla;